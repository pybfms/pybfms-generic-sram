/****************************************************************************
 * generic_sram_line_en_initiator_bfm.sv
 ****************************************************************************/

/**
 * Module: generic_sram_line_en_initiator_bfm
 * 
 * TODO: Add module documentation
 */
module generic_sram_line_en_initiator_bfm;


endmodule


